-- altera_cordic.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity altera_cordic is
	port (
		a      : in  std_logic_vector(15 downto 0) := (others => '0'); --      a.a
		areset : in  std_logic                     := '0';             -- areset.reset
		c      : out std_logic_vector(12 downto 0);                    --      c.c
		clk    : in  std_logic                     := '0';             --    clk.clk
		en     : in  std_logic_vector(0 downto 0)  := (others => '0'); --     en.en
		s      : out std_logic_vector(12 downto 0)                     --      s.s
	);
end entity altera_cordic;

architecture rtl of altera_cordic is
	component altera_cordic_CORDIC_0 is
		port (
			clk    : in  std_logic                     := 'X';             -- clk
			areset : in  std_logic                     := 'X';             -- reset
			en     : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- en
			a      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- a
			c      : out std_logic_vector(12 downto 0);                    -- c
			s      : out std_logic_vector(12 downto 0)                     -- s
		);
	end component altera_cordic_CORDIC_0;

begin

	cordic_0 : component altera_cordic_CORDIC_0
		port map (
			clk    => clk,    --    clk.clk
			areset => areset, -- areset.reset
			en     => en,     --     en.en
			a      => a,      --      a.a
			c      => c,      --      c.c
			s      => s       --      s.s
		);

end architecture rtl; -- of altera_cordic
